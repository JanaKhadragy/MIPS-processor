library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity Reg_file is
end Reg_file;

architecture Behavioral of Reg_file is

begin


end Behavioral;

